// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"
// CREATED		"Sun Oct 14 08:48:05 2018"

module AdderWithDisplay(
	SW,
	HEX2,
	HEX5,
	HEX7,
	LEDR
);


input wire	[8:0] SW;
output wire	[6:0] HEX2;
output wire	[6:0] HEX5;
output wire	[6:0] HEX7;
output wire	[17:17] LEDR;

wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_225;
wire	SYNTHESIZED_WIRE_226;
wire	SYNTHESIZED_WIRE_3;
wire	SYNTHESIZED_WIRE_227;
wire	SYNTHESIZED_WIRE_228;
wire	SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_229;
wire	SYNTHESIZED_WIRE_230;
wire	SYNTHESIZED_WIRE_13;
wire	SYNTHESIZED_WIRE_14;
wire	SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_231;
wire	SYNTHESIZED_WIRE_22;
wire	SYNTHESIZED_WIRE_23;
wire	SYNTHESIZED_WIRE_232;
wire	SYNTHESIZED_WIRE_26;
wire	SYNTHESIZED_WIRE_27;
wire	SYNTHESIZED_WIRE_28;
wire	SYNTHESIZED_WIRE_233;
wire	SYNTHESIZED_WIRE_234;
wire	SYNTHESIZED_WIRE_37;
wire	SYNTHESIZED_WIRE_38;
wire	SYNTHESIZED_WIRE_235;
wire	SYNTHESIZED_WIRE_46;
wire	SYNTHESIZED_WIRE_47;
wire	SYNTHESIZED_WIRE_48;
wire	SYNTHESIZED_WIRE_50;
wire	SYNTHESIZED_WIRE_51;
wire	SYNTHESIZED_WIRE_53;
wire	SYNTHESIZED_WIRE_54;
wire	SYNTHESIZED_WIRE_55;
wire	SYNTHESIZED_WIRE_59;
wire	SYNTHESIZED_WIRE_60;
wire	SYNTHESIZED_WIRE_236;
wire	SYNTHESIZED_WIRE_63;
wire	SYNTHESIZED_WIRE_64;
wire	SYNTHESIZED_WIRE_65;
wire	SYNTHESIZED_WIRE_67;
wire	SYNTHESIZED_WIRE_68;
wire	SYNTHESIZED_WIRE_237;
wire	SYNTHESIZED_WIRE_238;
wire	SYNTHESIZED_WIRE_239;
wire	SYNTHESIZED_WIRE_240;
wire	SYNTHESIZED_WIRE_241;
wire	SYNTHESIZED_WIRE_242;
wire	SYNTHESIZED_WIRE_75;
wire	SYNTHESIZED_WIRE_243;
wire	SYNTHESIZED_WIRE_244;
wire	SYNTHESIZED_WIRE_81;
wire	SYNTHESIZED_WIRE_85;
wire	SYNTHESIZED_WIRE_245;
wire	SYNTHESIZED_WIRE_95;
wire	SYNTHESIZED_WIRE_96;
wire	SYNTHESIZED_WIRE_97;
wire	SYNTHESIZED_WIRE_246;
wire	SYNTHESIZED_WIRE_107;
wire	SYNTHESIZED_WIRE_108;
wire	SYNTHESIZED_WIRE_247;
wire	SYNTHESIZED_WIRE_111;
wire	SYNTHESIZED_WIRE_112;
wire	SYNTHESIZED_WIRE_113;
wire	SYNTHESIZED_WIRE_248;
wire	SYNTHESIZED_WIRE_249;
wire	SYNTHESIZED_WIRE_129;
wire	SYNTHESIZED_WIRE_130;
wire	SYNTHESIZED_WIRE_250;
wire	SYNTHESIZED_WIRE_140;
wire	SYNTHESIZED_WIRE_251;
wire	SYNTHESIZED_WIRE_144;
wire	SYNTHESIZED_WIRE_145;
wire	SYNTHESIZED_WIRE_146;
wire	SYNTHESIZED_WIRE_147;
wire	SYNTHESIZED_WIRE_154;
wire	SYNTHESIZED_WIRE_155;
wire	SYNTHESIZED_WIRE_156;
wire	SYNTHESIZED_WIRE_159;
wire	SYNTHESIZED_WIRE_160;
wire	SYNTHESIZED_WIRE_161;
wire	SYNTHESIZED_WIRE_252;
wire	SYNTHESIZED_WIRE_253;
wire	SYNTHESIZED_WIRE_169;
wire	SYNTHESIZED_WIRE_254;
wire	SYNTHESIZED_WIRE_171;
wire	SYNTHESIZED_WIRE_172;
wire	SYNTHESIZED_WIRE_255;
wire	SYNTHESIZED_WIRE_174;
wire	SYNTHESIZED_WIRE_256;
wire	SYNTHESIZED_WIRE_180;
wire	SYNTHESIZED_WIRE_181;
wire	SYNTHESIZED_WIRE_182;
wire	SYNTHESIZED_WIRE_257;
wire	SYNTHESIZED_WIRE_189;
wire	SYNTHESIZED_WIRE_190;
wire	SYNTHESIZED_WIRE_191;
wire	SYNTHESIZED_WIRE_192;
wire	SYNTHESIZED_WIRE_258;
wire	SYNTHESIZED_WIRE_195;
wire	SYNTHESIZED_WIRE_196;
wire	SYNTHESIZED_WIRE_197;
wire	SYNTHESIZED_WIRE_259;
wire	SYNTHESIZED_WIRE_260;
wire	SYNTHESIZED_WIRE_205;
wire	SYNTHESIZED_WIRE_206;
wire	SYNTHESIZED_WIRE_261;
wire	SYNTHESIZED_WIRE_214;
wire	SYNTHESIZED_WIRE_215;
wire	SYNTHESIZED_WIRE_216;
wire	SYNTHESIZED_WIRE_219;
wire	SYNTHESIZED_WIRE_220;
wire	SYNTHESIZED_WIRE_221;




assign	SYNTHESIZED_WIRE_0 = SW[1] ^ SW[5];

assign	SYNTHESIZED_WIRE_237 = SYNTHESIZED_WIRE_0 ^ SW[0];

assign	SYNTHESIZED_WIRE_51 = SW[2] & SW[6];

assign	SYNTHESIZED_WIRE_225 =  ~SW[7];

assign	SYNTHESIZED_WIRE_227 =  ~SW[8];

assign	SYNTHESIZED_WIRE_6 = SYNTHESIZED_WIRE_225 & SYNTHESIZED_WIRE_226;

assign	HEX5[6] = SYNTHESIZED_WIRE_3 & SYNTHESIZED_WIRE_227;

assign	SYNTHESIZED_WIRE_228 = SW[7] & SW[6] & SW[5];

assign	SYNTHESIZED_WIRE_3 = SYNTHESIZED_WIRE_228 | SYNTHESIZED_WIRE_6;

assign	SYNTHESIZED_WIRE_231 = SW[8] & SW[7] & SYNTHESIZED_WIRE_226;

assign	SYNTHESIZED_WIRE_14 = SYNTHESIZED_WIRE_227 & SW[6] & SW[5];

assign	SYNTHESIZED_WIRE_230 = SYNTHESIZED_WIRE_227 & SYNTHESIZED_WIRE_225;

assign	SYNTHESIZED_WIRE_13 = SW[6] | SW[5];

assign	SYNTHESIZED_WIRE_50 = SW[2] & SYNTHESIZED_WIRE_229;

assign	SYNTHESIZED_WIRE_15 = SYNTHESIZED_WIRE_230 & SYNTHESIZED_WIRE_13;

assign	HEX5[5] = SYNTHESIZED_WIRE_14 | SYNTHESIZED_WIRE_15 | SYNTHESIZED_WIRE_231;

assign	SYNTHESIZED_WIRE_232 = SYNTHESIZED_WIRE_227 & SW[7] & SYNTHESIZED_WIRE_226;

assign	SYNTHESIZED_WIRE_22 = SYNTHESIZED_WIRE_225 & SYNTHESIZED_WIRE_226 & SW[5];

assign	SYNTHESIZED_WIRE_23 = SYNTHESIZED_WIRE_227 & SW[5];

assign	HEX5[4] = SYNTHESIZED_WIRE_22 | SYNTHESIZED_WIRE_23 | SYNTHESIZED_WIRE_232;

assign	HEX5[3] = SYNTHESIZED_WIRE_228 | SYNTHESIZED_WIRE_26 | SYNTHESIZED_WIRE_27;

assign	SYNTHESIZED_WIRE_26 = SYNTHESIZED_WIRE_28 & SYNTHESIZED_WIRE_233;

assign	SYNTHESIZED_WIRE_28 = SYNTHESIZED_WIRE_234 | SYNTHESIZED_WIRE_232;

assign	SYNTHESIZED_WIRE_234 = SW[8] & SYNTHESIZED_WIRE_225 & SW[6];

assign	SYNTHESIZED_WIRE_59 = SW[6] & SYNTHESIZED_WIRE_229;

assign	SYNTHESIZED_WIRE_235 = SW[8] & SW[7] & SYNTHESIZED_WIRE_233;

assign	SYNTHESIZED_WIRE_37 = SW[8] & SW[7] & SW[6];

assign	SYNTHESIZED_WIRE_38 = SYNTHESIZED_WIRE_230 & SW[6] & SYNTHESIZED_WIRE_233;

assign	HEX5[2] = SYNTHESIZED_WIRE_37 | SYNTHESIZED_WIRE_38 | SYNTHESIZED_WIRE_235;

assign	SYNTHESIZED_WIRE_55 = SW[7] & SW[6] & SYNTHESIZED_WIRE_233;

assign	SYNTHESIZED_WIRE_53 = SW[8] & SW[6] & SW[5];

assign	SYNTHESIZED_WIRE_54 = SYNTHESIZED_WIRE_232 & SW[5];

assign	SYNTHESIZED_WIRE_46 = SW[7] & SYNTHESIZED_WIRE_226 & SYNTHESIZED_WIRE_233;

assign	SYNTHESIZED_WIRE_47 = SYNTHESIZED_WIRE_230 & SYNTHESIZED_WIRE_226 & SW[5];

assign	HEX5[0] = SYNTHESIZED_WIRE_46 | SYNTHESIZED_WIRE_47 | SYNTHESIZED_WIRE_48 | SYNTHESIZED_WIRE_231;

assign	SYNTHESIZED_WIRE_60 = SYNTHESIZED_WIRE_50 | SYNTHESIZED_WIRE_51;

assign	HEX5[1] = SYNTHESIZED_WIRE_235 | SYNTHESIZED_WIRE_53 | SYNTHESIZED_WIRE_54 | SYNTHESIZED_WIRE_55;

assign	SYNTHESIZED_WIRE_48 = SYNTHESIZED_WIRE_234 & SW[5];

assign	SYNTHESIZED_WIRE_27 = SYNTHESIZED_WIRE_225 & SYNTHESIZED_WIRE_226 & SW[5];

assign	SYNTHESIZED_WIRE_236 = SYNTHESIZED_WIRE_59 | SYNTHESIZED_WIRE_60;

assign	SYNTHESIZED_WIRE_85 = SW[3] ^ SW[7];

assign	SYNTHESIZED_WIRE_64 = SW[3] & SW[7];

assign	SYNTHESIZED_WIRE_63 = SW[3] & SYNTHESIZED_WIRE_236;

assign	SYNTHESIZED_WIRE_67 = SW[7] & SYNTHESIZED_WIRE_236;

assign	SYNTHESIZED_WIRE_68 = SYNTHESIZED_WIRE_63 | SYNTHESIZED_WIRE_64;

assign	SYNTHESIZED_WIRE_238 = SYNTHESIZED_WIRE_65 ^ SYNTHESIZED_WIRE_229;

assign	SYNTHESIZED_WIRE_251 = SYNTHESIZED_WIRE_67 | SYNTHESIZED_WIRE_68;

assign	SYNTHESIZED_WIRE_248 =  ~SYNTHESIZED_WIRE_237;

assign	SYNTHESIZED_WIRE_242 =  ~SYNTHESIZED_WIRE_238;

assign	SYNTHESIZED_WIRE_241 =  ~SYNTHESIZED_WIRE_239;

assign	SYNTHESIZED_WIRE_243 =  ~SYNTHESIZED_WIRE_240;

assign	SYNTHESIZED_WIRE_81 = SYNTHESIZED_WIRE_241 & SYNTHESIZED_WIRE_242;

assign	HEX2[6] = SYNTHESIZED_WIRE_75 & SYNTHESIZED_WIRE_243;

assign	SYNTHESIZED_WIRE_244 = SYNTHESIZED_WIRE_239 & SYNTHESIZED_WIRE_238 & SYNTHESIZED_WIRE_237;

assign	SYNTHESIZED_WIRE_75 = SYNTHESIZED_WIRE_244 | SYNTHESIZED_WIRE_81;

assign	SYNTHESIZED_WIRE_246 = SYNTHESIZED_WIRE_240 & SYNTHESIZED_WIRE_239 & SYNTHESIZED_WIRE_242;

assign	SYNTHESIZED_WIRE_239 = SYNTHESIZED_WIRE_85 ^ SYNTHESIZED_WIRE_236;

assign	SYNTHESIZED_WIRE_96 = SYNTHESIZED_WIRE_243 & SYNTHESIZED_WIRE_238 & SYNTHESIZED_WIRE_237;

assign	SYNTHESIZED_WIRE_245 = SYNTHESIZED_WIRE_243 & SYNTHESIZED_WIRE_241;

assign	SYNTHESIZED_WIRE_95 = SYNTHESIZED_WIRE_238 | SYNTHESIZED_WIRE_237;

assign	SYNTHESIZED_WIRE_97 = SYNTHESIZED_WIRE_245 & SYNTHESIZED_WIRE_95;

assign	HEX2[5] = SYNTHESIZED_WIRE_96 | SYNTHESIZED_WIRE_97 | SYNTHESIZED_WIRE_246;

assign	SYNTHESIZED_WIRE_247 = SYNTHESIZED_WIRE_243 & SYNTHESIZED_WIRE_239 & SYNTHESIZED_WIRE_242;

assign	SYNTHESIZED_WIRE_107 = SYNTHESIZED_WIRE_241 & SYNTHESIZED_WIRE_242 & SYNTHESIZED_WIRE_237;

assign	SYNTHESIZED_WIRE_108 = SYNTHESIZED_WIRE_243 & SYNTHESIZED_WIRE_237;

assign	HEX2[4] = SYNTHESIZED_WIRE_107 | SYNTHESIZED_WIRE_108 | SYNTHESIZED_WIRE_247;

assign	HEX2[3] = SYNTHESIZED_WIRE_244 | SYNTHESIZED_WIRE_111 | SYNTHESIZED_WIRE_112;

assign	SYNTHESIZED_WIRE_172 = SW[1] & SW[5];

assign	SYNTHESIZED_WIRE_111 = SYNTHESIZED_WIRE_113 & SYNTHESIZED_WIRE_248;

assign	SYNTHESIZED_WIRE_113 = SYNTHESIZED_WIRE_249 | SYNTHESIZED_WIRE_247;

assign	SYNTHESIZED_WIRE_249 = SYNTHESIZED_WIRE_240 & SYNTHESIZED_WIRE_241 & SYNTHESIZED_WIRE_238;

assign	SYNTHESIZED_WIRE_250 = SYNTHESIZED_WIRE_240 & SYNTHESIZED_WIRE_239 & SYNTHESIZED_WIRE_248;

assign	SYNTHESIZED_WIRE_129 = SYNTHESIZED_WIRE_240 & SYNTHESIZED_WIRE_239 & SYNTHESIZED_WIRE_238;

assign	SYNTHESIZED_WIRE_130 = SYNTHESIZED_WIRE_245 & SYNTHESIZED_WIRE_238 & SYNTHESIZED_WIRE_248;

assign	HEX2[2] = SYNTHESIZED_WIRE_129 | SYNTHESIZED_WIRE_130 | SYNTHESIZED_WIRE_250;

assign	SYNTHESIZED_WIRE_161 = SYNTHESIZED_WIRE_239 & SYNTHESIZED_WIRE_238 & SYNTHESIZED_WIRE_248;

assign	SYNTHESIZED_WIRE_159 = SYNTHESIZED_WIRE_240 & SYNTHESIZED_WIRE_238 & SYNTHESIZED_WIRE_237;

assign	SYNTHESIZED_WIRE_160 = SYNTHESIZED_WIRE_247 & SYNTHESIZED_WIRE_237;

assign	SYNTHESIZED_WIRE_171 = SW[1] & SW[0];

assign	SYNTHESIZED_WIRE_140 = SW[4] ^ SW[8];

assign	SYNTHESIZED_WIRE_240 = SYNTHESIZED_WIRE_140 ^ SYNTHESIZED_WIRE_251;

assign	SYNTHESIZED_WIRE_145 = SW[4] & SW[8];

assign	SYNTHESIZED_WIRE_144 = SW[4] & SYNTHESIZED_WIRE_251;

assign	SYNTHESIZED_WIRE_146 = SW[8] & SYNTHESIZED_WIRE_251;

assign	SYNTHESIZED_WIRE_147 = SYNTHESIZED_WIRE_144 | SYNTHESIZED_WIRE_145;

assign	LEDR = SYNTHESIZED_WIRE_146 | SYNTHESIZED_WIRE_147;

assign	SYNTHESIZED_WIRE_154 = SYNTHESIZED_WIRE_239 & SYNTHESIZED_WIRE_242 & SYNTHESIZED_WIRE_248;

assign	SYNTHESIZED_WIRE_155 = SYNTHESIZED_WIRE_245 & SYNTHESIZED_WIRE_242 & SYNTHESIZED_WIRE_237;

assign	HEX2[0] = SYNTHESIZED_WIRE_154 | SYNTHESIZED_WIRE_155 | SYNTHESIZED_WIRE_156 | SYNTHESIZED_WIRE_246;

assign	SYNTHESIZED_WIRE_189 = SW[5] & SW[0];

assign	HEX2[1] = SYNTHESIZED_WIRE_250 | SYNTHESIZED_WIRE_159 | SYNTHESIZED_WIRE_160 | SYNTHESIZED_WIRE_161;

assign	SYNTHESIZED_WIRE_156 = SYNTHESIZED_WIRE_249 & SYNTHESIZED_WIRE_237;

assign	SYNTHESIZED_WIRE_112 = SYNTHESIZED_WIRE_241 & SYNTHESIZED_WIRE_242 & SYNTHESIZED_WIRE_237;

assign	SYNTHESIZED_WIRE_259 =  ~SW[1];

assign	SYNTHESIZED_WIRE_253 =  ~SW[2];

assign	SYNTHESIZED_WIRE_252 =  ~SW[3];

assign	SYNTHESIZED_WIRE_254 =  ~SW[4];

assign	SYNTHESIZED_WIRE_174 = SYNTHESIZED_WIRE_252 & SYNTHESIZED_WIRE_253;

assign	HEX7[6] = SYNTHESIZED_WIRE_169 & SYNTHESIZED_WIRE_254;

assign	SYNTHESIZED_WIRE_255 = SW[3] & SW[2] & SW[1];

assign	SYNTHESIZED_WIRE_190 = SYNTHESIZED_WIRE_171 | SYNTHESIZED_WIRE_172;

assign	SYNTHESIZED_WIRE_169 = SYNTHESIZED_WIRE_255 | SYNTHESIZED_WIRE_174;

assign	SYNTHESIZED_WIRE_257 = SW[4] & SW[3] & SYNTHESIZED_WIRE_253;

assign	SYNTHESIZED_WIRE_181 = SYNTHESIZED_WIRE_254 & SW[2] & SW[1];

assign	SYNTHESIZED_WIRE_256 = SYNTHESIZED_WIRE_254 & SYNTHESIZED_WIRE_252;

assign	SYNTHESIZED_WIRE_180 = SW[2] | SW[1];

assign	SYNTHESIZED_WIRE_182 = SYNTHESIZED_WIRE_256 & SYNTHESIZED_WIRE_180;

assign	HEX7[5] = SYNTHESIZED_WIRE_181 | SYNTHESIZED_WIRE_182 | SYNTHESIZED_WIRE_257;

assign	SYNTHESIZED_WIRE_258 = SYNTHESIZED_WIRE_254 & SW[3] & SYNTHESIZED_WIRE_253;

assign	SYNTHESIZED_WIRE_191 = SYNTHESIZED_WIRE_252 & SYNTHESIZED_WIRE_253 & SW[1];

assign	SYNTHESIZED_WIRE_192 = SYNTHESIZED_WIRE_254 & SW[1];

assign	SYNTHESIZED_WIRE_229 = SYNTHESIZED_WIRE_189 | SYNTHESIZED_WIRE_190;

assign	HEX7[4] = SYNTHESIZED_WIRE_191 | SYNTHESIZED_WIRE_192 | SYNTHESIZED_WIRE_258;

assign	HEX7[3] = SYNTHESIZED_WIRE_255 | SYNTHESIZED_WIRE_195 | SYNTHESIZED_WIRE_196;

assign	SYNTHESIZED_WIRE_195 = SYNTHESIZED_WIRE_197 & SYNTHESIZED_WIRE_259;

assign	SYNTHESIZED_WIRE_197 = SYNTHESIZED_WIRE_260 | SYNTHESIZED_WIRE_258;

assign	SYNTHESIZED_WIRE_260 = SW[4] & SYNTHESIZED_WIRE_252 & SW[2];

assign	SYNTHESIZED_WIRE_261 = SW[4] & SW[3] & SYNTHESIZED_WIRE_259;

assign	SYNTHESIZED_WIRE_205 = SW[4] & SW[3] & SW[2];

assign	SYNTHESIZED_WIRE_206 = SYNTHESIZED_WIRE_256 & SW[2] & SYNTHESIZED_WIRE_259;

assign	HEX7[2] = SYNTHESIZED_WIRE_205 | SYNTHESIZED_WIRE_206 | SYNTHESIZED_WIRE_261;

assign	SYNTHESIZED_WIRE_221 = SW[3] & SW[2] & SYNTHESIZED_WIRE_259;

assign	SYNTHESIZED_WIRE_65 = SW[2] ^ SW[6];

assign	SYNTHESIZED_WIRE_219 = SW[4] & SW[2] & SW[1];

assign	SYNTHESIZED_WIRE_220 = SYNTHESIZED_WIRE_258 & SW[1];

assign	SYNTHESIZED_WIRE_214 = SW[3] & SYNTHESIZED_WIRE_253 & SYNTHESIZED_WIRE_259;

assign	SYNTHESIZED_WIRE_215 = SYNTHESIZED_WIRE_256 & SYNTHESIZED_WIRE_253 & SW[1];

assign	HEX7[0] = SYNTHESIZED_WIRE_214 | SYNTHESIZED_WIRE_215 | SYNTHESIZED_WIRE_216 | SYNTHESIZED_WIRE_257;

assign	HEX7[1] = SYNTHESIZED_WIRE_261 | SYNTHESIZED_WIRE_219 | SYNTHESIZED_WIRE_220 | SYNTHESIZED_WIRE_221;

assign	SYNTHESIZED_WIRE_216 = SYNTHESIZED_WIRE_260 & SW[1];

assign	SYNTHESIZED_WIRE_196 = SYNTHESIZED_WIRE_252 & SYNTHESIZED_WIRE_253 & SW[1];

assign	SYNTHESIZED_WIRE_233 =  ~SW[5];

assign	SYNTHESIZED_WIRE_226 =  ~SW[6];


endmodule
