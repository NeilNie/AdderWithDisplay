// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"
// CREATED		"Wed Oct 10 11:07:41 2018"

module AdderWithDisplay(
	SW,
	HEX0
);


input wire	[6:0] SW;
output wire	[6:0] HEX0;

wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_79;
wire	SYNTHESIZED_WIRE_3;
wire	SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_5;
wire	SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_80;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_10;
wire	SYNTHESIZED_WIRE_11;
wire	SYNTHESIZED_WIRE_13;
wire	SYNTHESIZED_WIRE_14;
wire	SYNTHESIZED_WIRE_81;
wire	SYNTHESIZED_WIRE_82;
wire	SYNTHESIZED_WIRE_83;
wire	SYNTHESIZED_WIRE_84;
wire	SYNTHESIZED_WIRE_85;
wire	SYNTHESIZED_WIRE_21;
wire	SYNTHESIZED_WIRE_86;
wire	SYNTHESIZED_WIRE_87;
wire	SYNTHESIZED_WIRE_88;
wire	SYNTHESIZED_WIRE_89;
wire	SYNTHESIZED_WIRE_32;
wire	SYNTHESIZED_WIRE_33;
wire	SYNTHESIZED_WIRE_90;
wire	SYNTHESIZED_WIRE_91;
wire	SYNTHESIZED_WIRE_50;
wire	SYNTHESIZED_WIRE_55;
wire	SYNTHESIZED_WIRE_92;
wire	SYNTHESIZED_WIRE_62;
wire	SYNTHESIZED_WIRE_64;
wire	SYNTHESIZED_WIRE_65;
wire	SYNTHESIZED_WIRE_68;
wire	SYNTHESIZED_WIRE_69;
wire	SYNTHESIZED_WIRE_70;
wire	SYNTHESIZED_WIRE_71;
wire	SYNTHESIZED_WIRE_72;
wire	SYNTHESIZED_WIRE_73;
wire	SYNTHESIZED_WIRE_74;
wire	SYNTHESIZED_WIRE_75;
wire	SYNTHESIZED_WIRE_76;
wire	SYNTHESIZED_WIRE_77;
wire	SYNTHESIZED_WIRE_78;




assign	SYNTHESIZED_WIRE_0 = SW[1] ^ SW[2];

assign	SYNTHESIZED_WIRE_83 = SYNTHESIZED_WIRE_0 ^ SW[0];

assign	SYNTHESIZED_WIRE_4 = SW[3] & SW[4];

assign	SYNTHESIZED_WIRE_3 = SW[3] & SYNTHESIZED_WIRE_79;

assign	SYNTHESIZED_WIRE_5 = SW[4] & SYNTHESIZED_WIRE_79;

assign	SYNTHESIZED_WIRE_6 = SYNTHESIZED_WIRE_3 | SYNTHESIZED_WIRE_4;

assign	SYNTHESIZED_WIRE_80 = SYNTHESIZED_WIRE_5 | SYNTHESIZED_WIRE_6;

assign	SYNTHESIZED_WIRE_33 = SW[5] ^ SW[6];

assign	SYNTHESIZED_WIRE_10 = SW[5] & SW[6];

assign	SYNTHESIZED_WIRE_9 = SW[5] & SYNTHESIZED_WIRE_80;

assign	SYNTHESIZED_WIRE_13 = SW[6] & SYNTHESIZED_WIRE_80;

assign	SYNTHESIZED_WIRE_14 = SYNTHESIZED_WIRE_9 | SYNTHESIZED_WIRE_10;

assign	SYNTHESIZED_WIRE_81 = SYNTHESIZED_WIRE_11 ^ SYNTHESIZED_WIRE_79;

assign	SYNTHESIZED_WIRE_86 = SYNTHESIZED_WIRE_13 | SYNTHESIZED_WIRE_14;

assign	SYNTHESIZED_WIRE_88 =  ~SYNTHESIZED_WIRE_81;

assign	SYNTHESIZED_WIRE_84 =  ~SYNTHESIZED_WIRE_82;

assign	SYNTHESIZED_WIRE_21 = SYNTHESIZED_WIRE_82 & SYNTHESIZED_WIRE_83;

assign	SYNTHESIZED_WIRE_87 = SYNTHESIZED_WIRE_84 & SYNTHESIZED_WIRE_85;

assign	SYNTHESIZED_WIRE_68 = SYNTHESIZED_WIRE_21 | SYNTHESIZED_WIRE_81 | SYNTHESIZED_WIRE_86 | SYNTHESIZED_WIRE_87;

assign	SYNTHESIZED_WIRE_85 =  ~SYNTHESIZED_WIRE_83;

assign	SYNTHESIZED_WIRE_32 = SYNTHESIZED_WIRE_81 & SYNTHESIZED_WIRE_83;

assign	SYNTHESIZED_WIRE_89 = SYNTHESIZED_WIRE_88 & SYNTHESIZED_WIRE_85;

assign	SYNTHESIZED_WIRE_69 = SYNTHESIZED_WIRE_89 | SYNTHESIZED_WIRE_84 | SYNTHESIZED_WIRE_32;

assign	SYNTHESIZED_WIRE_82 = SYNTHESIZED_WIRE_33 ^ SYNTHESIZED_WIRE_80;

assign	SYNTHESIZED_WIRE_70 = SYNTHESIZED_WIRE_88 | SYNTHESIZED_WIRE_83 | SYNTHESIZED_WIRE_82;

assign	SYNTHESIZED_WIRE_90 = SYNTHESIZED_WIRE_81 & SYNTHESIZED_WIRE_85;

assign	SYNTHESIZED_WIRE_92 = SYNTHESIZED_WIRE_84 & SYNTHESIZED_WIRE_81;

assign	SYNTHESIZED_WIRE_62 = SYNTHESIZED_WIRE_83 & SYNTHESIZED_WIRE_88 & SYNTHESIZED_WIRE_82;

assign	SYNTHESIZED_WIRE_72 = SYNTHESIZED_WIRE_90 | SYNTHESIZED_WIRE_87;

assign	SYNTHESIZED_WIRE_73 = SYNTHESIZED_WIRE_89 | SYNTHESIZED_WIRE_91 | SYNTHESIZED_WIRE_86 | SYNTHESIZED_WIRE_50;

assign	SYNTHESIZED_WIRE_50 = SYNTHESIZED_WIRE_82 & SYNTHESIZED_WIRE_85;

assign	SYNTHESIZED_WIRE_91 = SYNTHESIZED_WIRE_82 & SYNTHESIZED_WIRE_88;

assign	SYNTHESIZED_WIRE_74 = SYNTHESIZED_WIRE_55 | SYNTHESIZED_WIRE_86 | SYNTHESIZED_WIRE_92 | SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_65 = SYNTHESIZED_WIRE_87 | SYNTHESIZED_WIRE_90 | SYNTHESIZED_WIRE_86;

assign	SYNTHESIZED_WIRE_76 = SW[1] & SW[2];

assign	SYNTHESIZED_WIRE_64 = SYNTHESIZED_WIRE_62 | SYNTHESIZED_WIRE_92;

assign	SYNTHESIZED_WIRE_71 = SYNTHESIZED_WIRE_64 | SYNTHESIZED_WIRE_65;

assign	SYNTHESIZED_WIRE_55 = SYNTHESIZED_WIRE_82 & SYNTHESIZED_WIRE_85;

assign	HEX0[0] =  ~SYNTHESIZED_WIRE_68;

assign	HEX0[1] =  ~SYNTHESIZED_WIRE_69;

assign	HEX0[2] =  ~SYNTHESIZED_WIRE_70;

assign	HEX0[3] =  ~SYNTHESIZED_WIRE_71;

assign	HEX0[4] =  ~SYNTHESIZED_WIRE_72;

assign	HEX0[5] =  ~SYNTHESIZED_WIRE_73;

assign	HEX0[6] =  ~SYNTHESIZED_WIRE_74;

assign	SYNTHESIZED_WIRE_75 = SW[1] & SW[0];

assign	SYNTHESIZED_WIRE_77 = SW[2] & SW[0];

assign	SYNTHESIZED_WIRE_78 = SYNTHESIZED_WIRE_75 | SYNTHESIZED_WIRE_76;

assign	SYNTHESIZED_WIRE_79 = SYNTHESIZED_WIRE_77 | SYNTHESIZED_WIRE_78;

assign	SYNTHESIZED_WIRE_11 = SW[3] ^ SW[4];


endmodule
